//`include "ALU_Decoder.sv"
//`include "Main_Decoder.sv"
//7
`timescale 1ns / 1ps
module Control_Unit_Top(Op,RegWrite,ImmSrc,ALUSrc,MemWrite,ResultSrc,Branch,funct3,funct7,ALUControl,PCSrc);

    input [6:0]Op,funct7;
    input [2:0]funct3;
    output RegWrite,ALUSrc,MemWrite,ResultSrc,Branch,PCSrc;
    output [1:0]ImmSrc;
    output [2:0]ALUControl;

    wire [1:0]ALUOp;

    Main_Decoder Main_Decoder(
                .Op(Op),
                .RegWrite(RegWrite),
                .ImmSrc(ImmSrc),
                .PCSrc(PCSrc),
                .MemWrite(MemWrite),
                .ResultSrc(ResultSrc),
                .Branch(Branch),
                .ALUSrc(ALUSrc),
                .ALUOp(ALUOp)
    );

    ALU_Decoder ALU_Decoder(
                            .ALUOp(ALUOp),
                            .funct3(funct3),
                            .funct7(funct7),
                            .op(Op),
                            .ALUControl(ALUControl)
    );


endmodule

////////////////////////////

module ALU_Decoder(ALUOp,funct3,funct7,op,ALUControl);

    input [1:0]ALUOp;
    input [2:0]funct3;
    input [6:0]funct7,op;
    output [2:0]ALUControl;

    wire cancatenation;
            
  assign cancatenation = {op,funct7};


assign ALUControl = (ALUOp == 2'b00) ? 3'b000 :
                    (ALUOp == 2'b01) ? 3'b001 :
                    ((ALUOp == 2'b10) & (funct3 == 3'b010)) ? 3'b101 :
                    ((ALUOp == 2'b10) & (funct3 == 3'b110)) ? 3'b011 :
                    ((ALUOp == 2'b10) & (funct3 == 3'b111)) ? 3'b010 :
                    ((ALUOp == 2'b10) & (funct3 == 3'b000) & (cancatenation == 2'b11)) ? 3'b001 :
                    /// here we not 11 the cancatenation to enable 00,01,10 //
                    ((ALUOp == 2'b10) & (funct3 == 3'b000) & (cancatenation != 2'b11)) ? 3'b000 : 3'b000;


    // Method 2
//    assign ALUControl = (ALUOp == 2'b00) ? 3'b000 :
//                        (ALUOp == 2'b01) ? 3'b001 :
//                        ((ALUOp == 2'b10) & (funct3 == 3'b000) & ({op[5],funct7[5]} == 2'b11)) ? 3'b001 : 
//                        ((ALUOp == 2'b10) & (funct3 == 3'b000) & ({op[5],funct7[5]} != 2'b11)) ? 3'b000 : 
//                        ((ALUOp == 2'b10) & (funct3 == 3'b010)) ? 3'b101 : 
//                        ((ALUOp == 2'b10) & (funct3 == 3'b110)) ? 3'b011 : 
//                        ((ALUOp == 2'b10) & (funct3 == 3'b111)) ? 3'b010 : 
//                                                                  3'b000 ;
endmodule

/////////////////////

module Main_Decoder(Op,RegWrite,ImmSrc,ALUSrc,MemWrite,ResultSrc,Branch,ALUOp, PCSrc);
    input [6:0]Op;
    output RegWrite,ALUSrc,MemWrite,ResultSrc,Branch, PCSrc;
    output [1:0]ImmSrc,ALUOp;
    
    assign PCSrc = Branch;
    
    assign RegWrite = (Op == 7'b0000011 | Op == 7'b0110011) ? 1'b1 :
                                                              1'b0 ;
    assign ImmSrc = (Op == 7'b0100011) ? 2'b01 : 
                    (Op == 7'b1100011) ? 2'b10 :    
                                         2'b00 ;
    assign ALUSrc = (Op == 7'b0000011 | Op == 7'b0100011) ? 1'b1 :
                                                            1'b0 ;
    assign MemWrite = (Op == 7'b0100011) ? 1'b1 :
                                           1'b0 ;
    assign ResultSrc = (Op == 7'b0000011) ? 1'b1 :
                                            1'b0 ;
    assign Branch = (Op == 7'b1100011) ? 1'b1 :
                                         1'b0 ;
    assign ALUOp = (Op == 7'b0110011) ? 2'b10 :
                   (Op == 7'b1100011) ? 2'b01 :
                                        2'b00 ;

endmodule